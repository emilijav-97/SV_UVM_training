interface inter_f(input logic clk, rst);
  
  bit valid_in;
  bit mem_full;
  
endinterface: inter_f