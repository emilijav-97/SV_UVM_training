module memory_driver
    (
      input clk,
      input rst,
      input valid_in,
      output mem_full
    );

endmodule